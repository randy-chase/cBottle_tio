netcdf file {
dimensions:
	pix = 49152 ;
	time = UNLIMITED ; // (40 currently)
	crs = 1 ;
variables:
	float crs(crs) ;
		crs:grid_mapping_name = "healpix" ;
		crs:healpix_nside = 64LL ;
		crs:healpix_order = "ring" ;
	int64 time(time) ;
		time:units = "seconds since 1970-1-1 0:0:0" ;
		time:calendar = "standard" ;
	float U1000(time, pix) ;
		U1000:_FillValue = NaNf ;
		U1000:grid_mapping = "crs" ;
	float U850(time, pix) ;
		U850:_FillValue = NaNf ;
		U850:grid_mapping = "crs" ;
	float U700(time, pix) ;
		U700:_FillValue = NaNf ;
		U700:grid_mapping = "crs" ;
	float U500(time, pix) ;
		U500:_FillValue = NaNf ;
		U500:grid_mapping = "crs" ;
	float U300(time, pix) ;
		U300:_FillValue = NaNf ;
		U300:grid_mapping = "crs" ;
	float U200(time, pix) ;
		U200:_FillValue = NaNf ;
		U200:grid_mapping = "crs" ;
	float U50(time, pix) ;
		U50:_FillValue = NaNf ;
		U50:grid_mapping = "crs" ;
	float U10(time, pix) ;
		U10:_FillValue = NaNf ;
		U10:grid_mapping = "crs" ;
	float V1000(time, pix) ;
		V1000:_FillValue = NaNf ;
		V1000:grid_mapping = "crs" ;
	float V850(time, pix) ;
		V850:_FillValue = NaNf ;
		V850:grid_mapping = "crs" ;
	float V700(time, pix) ;
		V700:_FillValue = NaNf ;
		V700:grid_mapping = "crs" ;
	float V500(time, pix) ;
		V500:_FillValue = NaNf ;
		V500:grid_mapping = "crs" ;
	float V300(time, pix) ;
		V300:_FillValue = NaNf ;
		V300:grid_mapping = "crs" ;
	float V200(time, pix) ;
		V200:_FillValue = NaNf ;
		V200:grid_mapping = "crs" ;
	float V50(time, pix) ;
		V50:_FillValue = NaNf ;
		V50:grid_mapping = "crs" ;
	float V10(time, pix) ;
		V10:_FillValue = NaNf ;
		V10:grid_mapping = "crs" ;
	float T1000(time, pix) ;
		T1000:_FillValue = NaNf ;
		T1000:grid_mapping = "crs" ;
	float T850(time, pix) ;
		T850:_FillValue = NaNf ;
		T850:grid_mapping = "crs" ;
	float T700(time, pix) ;
		T700:_FillValue = NaNf ;
		T700:grid_mapping = "crs" ;
	float T500(time, pix) ;
		T500:_FillValue = NaNf ;
		T500:grid_mapping = "crs" ;
	float T300(time, pix) ;
		T300:_FillValue = NaNf ;
		T300:grid_mapping = "crs" ;
	float T200(time, pix) ;
		T200:_FillValue = NaNf ;
		T200:grid_mapping = "crs" ;
	float T50(time, pix) ;
		T50:_FillValue = NaNf ;
		T50:grid_mapping = "crs" ;
	float T10(time, pix) ;
		T10:_FillValue = NaNf ;
		T10:grid_mapping = "crs" ;
	float Z1000(time, pix) ;
		Z1000:_FillValue = NaNf ;
		Z1000:grid_mapping = "crs" ;
	float Z850(time, pix) ;
		Z850:_FillValue = NaNf ;
		Z850:grid_mapping = "crs" ;
	float Z700(time, pix) ;
		Z700:_FillValue = NaNf ;
		Z700:grid_mapping = "crs" ;
	float Z500(time, pix) ;
		Z500:_FillValue = NaNf ;
		Z500:grid_mapping = "crs" ;
	float Z300(time, pix) ;
		Z300:_FillValue = NaNf ;
		Z300:grid_mapping = "crs" ;
	float Z200(time, pix) ;
		Z200:_FillValue = NaNf ;
		Z200:grid_mapping = "crs" ;
	float Z50(time, pix) ;
		Z50:_FillValue = NaNf ;
		Z50:grid_mapping = "crs" ;
	float Z10(time, pix) ;
		Z10:_FillValue = NaNf ;
		Z10:grid_mapping = "crs" ;
	float tcwv(time, pix) ;
		tcwv:_FillValue = NaNf ;
		tcwv:grid_mapping = "crs" ;
	float cllvi(time, pix) ;
		cllvi:_FillValue = NaNf ;
		cllvi:grid_mapping = "crs" ;
	float clivi(time, pix) ;
		clivi:_FillValue = NaNf ;
		clivi:grid_mapping = "crs" ;
	float tas(time, pix) ;
		tas:_FillValue = NaNf ;
		tas:grid_mapping = "crs" ;
	float uas(time, pix) ;
		uas:_FillValue = NaNf ;
		uas:grid_mapping = "crs" ;
	float vas(time, pix) ;
		vas:_FillValue = NaNf ;
		vas:grid_mapping = "crs" ;
	float rlut(time, pix) ;
		rlut:_FillValue = NaNf ;
		rlut:grid_mapping = "crs" ;
	float rsut(time, pix) ;
		rsut:_FillValue = NaNf ;
		rsut:grid_mapping = "crs" ;
	float pres_msl(time, pix) ;
		pres_msl:_FillValue = NaNf ;
		pres_msl:grid_mapping = "crs" ;
	float pr(time, pix) ;
		pr:_FillValue = NaNf ;
		pr:grid_mapping = "crs" ;
	float rsds(time, pix) ;
		rsds:_FillValue = NaNf ;
		rsds:grid_mapping = "crs" ;
	float sst(time, pix) ;
		sst:_FillValue = NaNf ;
		sst:grid_mapping = "crs" ;
	float sic(time, pix) ;
		sic:_FillValue = NaNf ;
		sic:grid_mapping = "crs" ;

// global attributes:
		:history = "scripts/inference_coarse.py /tmp/out.cbottle --dataset amip /tmp/amip/ --sample.batch_gpu 4 --sample.seed 0 --sample.bf16 --sample.sigma_max 1000" ;
data:
	time = 0, 1, 2, 3;
}
